module binding_module;
bind aes_binary v_aes_binary s_aes_binary( clk, data_stable, key_ready, finished,round_type_sel);  
endmodule
