module binding_module;
bind RSA_binary v_RSA_binary s_RSA_binary( clk, data_stable,	key_ready, finished,round_type_sel);  
endmodule
